`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   06:59:05 10/22/2022
// Design Name:   mux64_32
// Module Name:   E:/University/computer_architecture_lab/mips/test.v
// Project Name:  mips
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: mux64_32
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////
`include "mux64_32.v"
module mux_test;

	// Inputs
	reg [31:0] a;
	reg [31:0] b;
	reg s;

	// Outputs
	wire [31:0] c;

	// Instantiate the Unit Under Test (UUT)
		initial begin
		$dumpfile("mux_test.vcd");
		$dumpvars(0, mux_test);
	end
	mux64_32 uut (
		.a(a), 
		.b(b), 
		.s(s), 
		.c(c)
	);

	initial begin
		// Initialize Inputs
		a = 0;
		b = 40;
		s = 1;

		// Wait 100 ns for global reset to finish
		#100;
        
		a = 30;
		b = 0;
		s = 0;

		// Wait 100 ns for global reset to finish
		#100;

	end
      
endmodule

